�PNG

   IHDR  ,   #   .\7   	pHYs  M  uQJ��   tEXtSoftware Adobe ImageReadyq�e<  FIDATx���1o�@��bÖ�:�Tl�4�R$6Č�H2�T���Kg$6� �1�H����tB�[%��XN�/Vb�I��Mq��I|w�ދ                      ,�E���{7ѿ����z����~��ı�P���W���:��X;�6���V=����ۧ��^�BU��)�ud���B����AbbS�9Ff��2� ,��?��f;9�te���a8�<��������ݳ	q�����u>~H��v/�/�BZω
&EY�LӢ
��e{q�	��몟�9�ӝ���J-���d[���/����_�?����z� n��!0����6	�7�כ-y�j�7pݴ��ū���a ��
��m��~�����V��b�Q6KG��9��H�(k8<�Ǝa��l���|�rp�]������4L�t�ϖ��,	MlĖ�-%\=�A˺�5/��Y��b���D�Z�3T���*<���`:Ң��}M:�DE
A�au�i��l[����7��f'-�`��F~|������0J�O�����ͦ���WDʬ!;}�                  ���~�uI6S�    IEND�B`�